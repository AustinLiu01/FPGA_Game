module Display_double(in, out);
	input [5:0]in ;
	output reg [13:0]out;
	
	always @(*) begin
		case(in)
			6'b000000: out = {7'b1000000 , 7'b1000000 } ;
			6'b000001: out = {7'b1000000 , 7'b1111001 } ;
			6'b000010: out = {7'b1000000 , 7'b0100100 } ;
			6'b000011: out = {7'b1000000 , 7'b0110000 } ;
			6'b000100: out = {7'b1000000 , 7'b0011001 } ;
			6'b000101: out = {7'b1000000 , 7'b0010010 } ;
			6'b000110: out = {7'b1000000 , 7'b0000010 } ;
			6'b000111: out = {7'b1000000 , 7'b1111000 } ;
			6'b001000: out = {7'b1000000 , 7'b0000000 } ;
			6'b001001: out = {7'b1000000 , 7'b0010000 } ;
			6'b001010: out = {7'b1111001 , 7'b1000000 } ;
			6'b001011: out = {7'b1111001 , 7'b1111001 } ;
			6'b001100: out = {7'b1111001 , 7'b0100100 } ;
			6'b001101: out = {7'b1111001 , 7'b0110000 } ;
			6'b001110: out = {7'b1111001 , 7'b0011001 } ;
			6'b001111: out = {7'b1111001 , 7'b0010010 } ;
			6'b010000: out = {7'b1111001 , 7'b0000010 } ;
			6'b010001: out = {7'b1111001 , 7'b1111000 } ;
			6'b010010: out = {7'b1111001 , 7'b0000000 } ;
			6'b010011: out = {7'b1111001 , 7'b0010000 } ;
			6'b010100: out = {7'b0100100 , 7'b1000000 } ;
			6'b010101: out = {7'b0100100 , 7'b1111001 } ;
			6'b010110: out = {7'b0100100 , 7'b0100100 } ;
			6'b010111: out = {7'b0100100 , 7'b0110000 } ;
			6'b011000: out = {7'b0100100 , 7'b0011001 } ;
			6'b011001: out = {7'b0100100 , 7'b0010010 } ;
			6'b011010: out = {7'b0100100 , 7'b0000010 } ;
			6'b011011: out = {7'b0100100 , 7'b1111000 } ;
			6'b011100: out = {7'b0100100 , 7'b0000000 } ;
			6'b011101: out = {7'b0100100 , 7'b0010000 } ;
			6'b011110: out = {7'b0110000 , 7'b1000000 } ;
			6'b011111: out = {7'b0110000 , 7'b1111001 } ;
			6'b100000: out = {7'b0110000 , 7'b0100100 } ;
			6'b100001: out = {7'b0110000 , 7'b0110000 } ;
			6'b100010: out = {7'b0110000 , 7'b0011001 } ;
			6'b100011: out = {7'b0110000 , 7'b0010010 } ;
			6'b100100: out = {7'b0110000 , 7'b0000010 } ;
			6'b100101: out = {7'b0110000 , 7'b1111000 } ;
			6'b100110: out = {7'b0110000 , 7'b0000000 } ;
			6'b100111: out = {7'b0110000 , 7'b0010000 } ;
			6'b101000: out = {7'b0011001 , 7'b1000000 } ;
			6'b101001: out = {7'b0011001 , 7'b1111001 } ;
			6'b101010: out = {7'b0011001 , 7'b0100100 } ;
			6'b101011: out = {7'b0011001 , 7'b0110000 } ;
			6'b101100: out = {7'b0011001 , 7'b0011001 } ;
			6'b101101: out = {7'b0011001 , 7'b0010010 } ;
			6'b101110: out = {7'b0011001 , 7'b0000010 } ;
			6'b101111: out = {7'b0011001 , 7'b1111000 } ;
			6'b110000: out = {7'b0011001 , 7'b0000000 } ;
			6'b110001: out = {7'b0011001 , 7'b0010000 } ;
			6'b110010: out = {7'b0010010 , 7'b1000000 } ;
		endcase
	end
endmodule
