module Sum_10(in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, sum);
	input [5:0]in_0;
	input [5:0]in_1;
	input [5:0]in_2;
	input [5:0]in_3;
	input [5:0]in_4;
	input [5:0]in_5;
	input [5:0]in_6;
	input [5:0]in_7;
	input [5:0]in_8;
	input [5:0]in_9;
	
	output [5:0]sum;
	
	assign sum = in_0 + in_1 +in_2 + in_3 + in_4 + in_5 + in_6 + in_7 + in_8 + in_9 ;
	
	

endmodule
